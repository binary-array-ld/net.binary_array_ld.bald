netcdf ogcClassC {
dimensions:
        d0 = 1 ;
	d1 = 1 ;
variables:
	int var0 ;
	int var1 ;
:title = "Sample netCDF file definition with alias terms from the netCDF user guide" ;
data:
}
