netcdf attributes {
    dimensions:
        d0 = 10 ;
        d1 = 90 ;
        d2 = 15 ;
        d3 = 60 ;
    variables:
        int var0(d0, d1, d2) ;
            var0:test__references = "var1 var2" ;
            var0:test__name = "var0" ;
        int var1(d1, d2, d3) ;
            var1:test__references = "var2";
        int var2(d2) ;

    :bald__isPrefixedBy = "prefix_list";

    group: prefix_list {
        :bald__ = "https://www.opengis.net/def/binary-array-ld/";
        :test__ = "http://test.binary-array-ld.net/vocab/";
    }
}